library verilog;
use verilog.vl_types.all;
entity channel_sel is
    generic(
        MAX_SYNC_NUM    : integer := 26;
        ch1_addr_base   : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch2_addr_base   : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch3_addr_base   : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch4_addr_base   : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch5_addr_base   : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch6_addr_base   : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch7_addr_base   : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch8_addr_base   : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch9_addr_base   : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch10_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch11_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch12_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch13_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch14_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch15_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch16_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch17_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch18_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch19_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch20_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch21_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch22_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch23_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch24_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ch25_addr_base  : vl_logic_vector(0 to 19) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0)
    );
    port(
        clk             : in     vl_logic;
        ch_sgn_in       : in     vl_logic_vector(14 downto 0);
        ch_sgn_out      : out    vl_logic;
        ch_sync_in      : in     vl_logic;
        ch_c_in         : in     vl_logic_vector(2 downto 0);
        ch_sync_out     : out    vl_logic;
        mcu_n_rst       : in     vl_logic;
        mcu_data        : out    vl_logic_vector(7 downto 0);
        mcu_start       : in     vl_logic;
        mcu_end         : out    vl_logic;
        mcu_data_sel    : in     vl_logic_vector(2 downto 0);
        addr_base       : out    vl_logic_vector(19 downto 0);
        mem_data        : in     vl_logic_vector(7 downto 0);
        sample_en       : out    vl_logic;
        pulse_cnt       : in     vl_logic_vector(15 downto 0);
        sync_cnt_out    : out    vl_logic_vector(7 downto 0);
        clk_cnt         : in     vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of MAX_SYNC_NUM : constant is 1;
    attribute mti_svvh_generic_type of ch1_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch2_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch3_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch4_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch5_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch6_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch7_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch8_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch9_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch10_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch11_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch12_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch13_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch14_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch15_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch16_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch17_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch18_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch19_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch20_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch21_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch22_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch23_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch24_addr_base : constant is 1;
    attribute mti_svvh_generic_type of ch25_addr_base : constant is 1;
end channel_sel;
