library verilog;
use verilog.vl_types.all;
entity maxii_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end maxii_routing_wire;
